// opcodes.svh

/*
Contains typedef for top-level operations
*/

`ifndef _OPCODES_SVH_
`define _OPCODES_SVH_

typedef enum {
    ADD,
    SUB,
    MUL,
    DIV
} opcodes;

`endif  // _OPCODES_SVH_
